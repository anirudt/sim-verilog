module comp4(a,b,g,e,l);
	input [3:0] a,b;
	output reg g,e,l;

	initial begin g<=0;e=1;l=0; end

	